`define HADDR_SIZE 32
`define HDATA_SIZE 32
`define PADDR_SIZE 10
`define PDATA_SIZE  8
`define SYNC_DEPTH  3